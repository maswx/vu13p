// create by 小火车(masw@masw.tech)
//
module xdma_ddr4x4_top (
  output           c0_ddr4_act_n   ,
  output   [16:0]  c0_ddr4_adr     ,
  output   [ 1:0]  c0_ddr4_ba      ,
  output   [ 0:0]  c0_ddr4_bg      ,
  output   [ 0:0]  c0_ddr4_ck_c    ,
  output   [ 0:0]  c0_ddr4_ck_t    ,
  output   [ 0:0]  c0_ddr4_cke     ,
  input            c0_ddr4_clk_n   ,
  input            c0_ddr4_clk_p   ,
  output   [ 0:0]  c0_ddr4_cs_n    ,
  inout    [ 7:0]  c0_ddr4_dm_n    ,
  inout    [63:0]  c0_ddr4_dq      ,
  inout    [ 7:0]  c0_ddr4_dqs_c   ,
  inout    [ 7:0]  c0_ddr4_dqs_t   ,
  output   [ 0:0]  c0_ddr4_odt     ,
  output           c0_ddr4_reset_n ,

  output           c1_ddr4_act_n   ,
  output   [16:0]  c1_ddr4_adr     ,
  output   [ 1:0]  c1_ddr4_ba      ,
  output   [ 0:0]  c1_ddr4_bg      ,
  output   [ 0:0]  c1_ddr4_ck_c    ,
  output   [ 0:0]  c1_ddr4_ck_t    ,
  output   [ 0:0]  c1_ddr4_cke     ,
  input            c1_ddr4_clk_n   ,
  input            c1_ddr4_clk_p   ,
  output   [ 0:0]  c1_ddr4_cs_n    ,
  inout    [ 7:0]  c1_ddr4_dm_n    ,
  inout    [63:0]  c1_ddr4_dq      ,
  inout    [ 7:0]  c1_ddr4_dqs_c   ,
  inout    [ 7:0]  c1_ddr4_dqs_t   ,
  output   [ 0:0]  c1_ddr4_odt     ,
  output           c1_ddr4_reset_n ,

  output           c2_ddr4_act_n   ,
  output   [16:0]  c2_ddr4_adr     ,
  output   [ 1:0]  c2_ddr4_ba      ,
  output   [ 0:0]  c2_ddr4_bg      ,
  output   [ 0:0]  c2_ddr4_ck_c    ,
  output   [ 0:0]  c2_ddr4_ck_t    ,
  output   [ 0:0]  c2_ddr4_cke     ,
  input            c2_ddr4_clk_n   ,
  input            c2_ddr4_clk_p   ,
  output   [ 0:0]  c2_ddr4_cs_n    ,
  inout    [ 7:0]  c2_ddr4_dm_n    ,
  inout    [63:0]  c2_ddr4_dq      ,
  inout    [ 7:0]  c2_ddr4_dqs_c   ,
  inout    [ 7:0]  c2_ddr4_dqs_t   ,
  output   [ 0:0]  c2_ddr4_odt     ,
  output           c2_ddr4_reset_n ,

  output           c3_ddr4_act_n   ,
  output   [16:0]  c3_ddr4_adr     ,
  output   [ 1:0]  c3_ddr4_ba      ,
  output   [ 0:0]  c3_ddr4_bg      ,
  output   [ 0:0]  c3_ddr4_ck_c    ,
  output   [ 0:0]  c3_ddr4_ck_t    ,
  output   [ 0:0]  c3_ddr4_cke     ,
  input            c3_ddr4_clk_n   ,
  input            c3_ddr4_clk_p   ,
  output   [ 0:0]  c3_ddr4_cs_n    ,
  inout    [ 7:0]  c3_ddr4_dm_n    ,
  inout    [63:0]  c3_ddr4_dq      ,
  inout    [ 7:0]  c3_ddr4_dqs_c   ,
  inout    [ 7:0]  c3_ddr4_dqs_t   ,
  output   [ 0:0]  c3_ddr4_odt     ,
  output           c3_ddr4_reset_n ,


  input    [15:0]  pcie_lane_rxn   ,
  input    [15:0]  pcie_lane_rxp   ,
  output   [15:0]  pcie_lane_txn   ,
  output   [15:0]  pcie_lane_txp   ,
  input            pcie_perst_n    ,
  input    [ 0:0]  pcie_ref_clk_n  ,
  input    [ 0:0]  pcie_ref_clk_p  ,
  output           pcie_link_up    
);


//log by masw@masw.tech : 可以直接调用BD文件
xdma_ddr4x4 xdma_ddr4x4_i (
	.c0_ddr4_act_n        (c0_ddr4_act_n         ),
	.c0_ddr4_adr          (c0_ddr4_adr           ),
	.c0_ddr4_ba           (c0_ddr4_ba            ),
	.c0_ddr4_bg           (c0_ddr4_bg            ),
	.c0_ddr4_ck_c         (c0_ddr4_ck_c          ),
	.c0_ddr4_ck_t         (c0_ddr4_ck_t          ),
	.c0_ddr4_cke          (c0_ddr4_cke           ),
	.c0_ddr4_clk_clk_n    (c0_ddr4_clk_n         ),
	.c0_ddr4_clk_clk_p    (c0_ddr4_clk_p         ),
	.c0_ddr4_cs_n         (c0_ddr4_cs_n          ),
	.c0_ddr4_dm_n         (c0_ddr4_dm_n          ),
	.c0_ddr4_dq           (c0_ddr4_dq            ),
	.c0_ddr4_dqs_c        (c0_ddr4_dqs_c         ),
	.c0_ddr4_dqs_t        (c0_ddr4_dqs_t         ),
	.c0_ddr4_odt          (c0_ddr4_odt           ),
	.c0_ddr4_reset_n      (c0_ddr4_reset_n       ),
	.c1_ddr4_act_n        (c1_ddr4_act_n         ),
	.c1_ddr4_adr          (c1_ddr4_adr           ),
	.c1_ddr4_ba           (c1_ddr4_ba            ),
	.c1_ddr4_bg           (c1_ddr4_bg            ),
	.c1_ddr4_ck_c         (c1_ddr4_ck_c          ),
	.c1_ddr4_ck_t         (c1_ddr4_ck_t          ),
	.c1_ddr4_cke          (c1_ddr4_cke           ),
	.c1_ddr4_clk_clk_n    (c1_ddr4_clk_n         ),
	.c1_ddr4_clk_clk_p    (c1_ddr4_clk_p         ),
	.c1_ddr4_cs_n         (c1_ddr4_cs_n          ),
	.c1_ddr4_dm_n         (c1_ddr4_dm_n          ),
	.c1_ddr4_dq           (c1_ddr4_dq            ),
	.c1_ddr4_dqs_c        (c1_ddr4_dqs_c         ),
	.c1_ddr4_dqs_t        (c1_ddr4_dqs_t         ),
	.c1_ddr4_odt          (c1_ddr4_odt           ),
	.c1_ddr4_reset_n      (c1_ddr4_reset_n       ),
	.c2_ddr4_act_n        (c2_ddr4_act_n         ),
	.c2_ddr4_adr          (c2_ddr4_adr           ),
	.c2_ddr4_ba           (c2_ddr4_ba            ),
	.c2_ddr4_bg           (c2_ddr4_bg            ),
	.c2_ddr4_ck_c         (c2_ddr4_ck_c          ),
	.c2_ddr4_ck_t         (c2_ddr4_ck_t          ),
	.c2_ddr4_cke          (c2_ddr4_cke           ),
	.c2_ddr4_clk_clk_n    (c2_ddr4_clk_n         ),
	.c2_ddr4_clk_clk_p    (c2_ddr4_clk_p         ),
	.c2_ddr4_cs_n         (c2_ddr4_cs_n          ),
	.c2_ddr4_dm_n         (c2_ddr4_dm_n          ),
	.c2_ddr4_dq           (c2_ddr4_dq            ),
	.c2_ddr4_dqs_c        (c2_ddr4_dqs_c         ),
	.c2_ddr4_dqs_t        (c2_ddr4_dqs_t         ),
	.c2_ddr4_odt          (c2_ddr4_odt           ),
	.c2_ddr4_reset_n      (c2_ddr4_reset_n       ),
	.c3_ddr4_act_n        (c3_ddr4_act_n         ),
	.c3_ddr4_adr          (c3_ddr4_adr           ),
	.c3_ddr4_ba           (c3_ddr4_ba            ),
	.c3_ddr4_bg           (c3_ddr4_bg            ),
	.c3_ddr4_ck_c         (c3_ddr4_ck_c          ),
	.c3_ddr4_ck_t         (c3_ddr4_ck_t          ),
	.c3_ddr4_cke          (c3_ddr4_cke           ),
	.c3_ddr4_clk_clk_n    (c3_ddr4_clk_n         ),
	.c3_ddr4_clk_clk_p    (c3_ddr4_clk_p         ),
	.c3_ddr4_cs_n         (c3_ddr4_cs_n          ),
	.c3_ddr4_dm_n         (c3_ddr4_dm_n          ),
	.c3_ddr4_dq           (c3_ddr4_dq            ),
	.c3_ddr4_dqs_c        (c3_ddr4_dqs_c         ),
	.c3_ddr4_dqs_t        (c3_ddr4_dqs_t         ),
	.c3_ddr4_odt          (c3_ddr4_odt           ),
	.c3_ddr4_reset_n      (c3_ddr4_reset_n       ),
	.pcie_lane_rxn        (pcie_lane_rxn         ),
	.pcie_lane_rxp        (pcie_lane_rxp         ),
	.pcie_lane_txn        (pcie_lane_txn         ),
	.pcie_lane_txp        (pcie_lane_txp         ),
	.pcie_link_up         (pcie_link_up          ),
	.pcie_perst_n         (pcie_perst_n          ),
	.pcie_ref_clk_n       (pcie_ref_clk_n        ),
	.pcie_ref_clk_p       (pcie_ref_clk_p        )
);
endmodule
